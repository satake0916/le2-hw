library verilog;
use verilog.vl_types.all;
entity junjo_vlg_tst is
end junjo_vlg_tst;
