library verilog;
use verilog.vl_types.all;
entity fulladder_vlg_tst is
end fulladder_vlg_tst;
